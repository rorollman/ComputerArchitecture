module nor_1b(output C, input A, B);
	nor(C, A, B);
endmodule
