module not_1b(output B, input A);
	not(B, A);
endmodule
